module enc8to3(
    input [7:0]a,
    input en,
    output reg [2:0]y
);
always @(*)begin
    if(en)begin
        case(a)
        8'b00000000:y=3'b000;
        8'b00000001:y=3'b001;
        8'b00000010:y=3'b010;
        8'b00000011:y=3'b011;
        8'b00000100:y=3'b100;
        8'b00000101:y=3'b101; 
        8'b00000110:y=3'b110;
        8'b00000111:y=3'b111;
        default:y=3'b111;
        endcase
    end
    else
    begin
        y=3'b000;
    end
end
endmodule
