module par_mux_tb;
 parameter n=8;
 parameter m=3;

reg [7:0]in;
reg [2:0]sel;
wire y;

par_mux#(8) DUT(.*);

initial begin
$monitor ("$time=%0t  | in=%b sel=%b | y=%b",
$time,in,sel,y);
$dumpfile("par_mux.vcd");
$dumpvars(0,par_mux_tb);

in =8'b10001010;
sel = 3'b000; #10;
sel = 3'b001; #10;

in =8'b11001010;
sel = 3'b010; #10;
sel = 3'b011; #10;
sel = 3'b010; #10;
$finish;

end
endmodule
